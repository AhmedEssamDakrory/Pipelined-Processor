library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.Numeric_Std.all;
package Common is   
   type state_type is (st,wt,snt,wnt);
end Common;
package body Common is
end Common;